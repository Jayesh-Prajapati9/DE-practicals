<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-35.0062,-0.221008,182.84,-107.898</PageViewport>
<gate>
<ID>387</ID>
<type>GA_LED</type>
<position>50,-76.5</position>
<input>
<ID>N_in1</ID>154 </input>
<input>
<ID>N_in2</ID>154 </input>
<input>
<ID>N_in3</ID>154 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>-167.5,-45.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>AA_LABEL</type>
<position>-137,-46.5</position>
<gparam>LABEL_TEXT A'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>389</ID>
<type>GA_LED</type>
<position>50,-85</position>
<input>
<ID>N_in0</ID>153 </input>
<input>
<ID>N_in3</ID>153 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>390</ID>
<type>AA_LABEL</type>
<position>138.5,-12</position>
<gparam>LABEL_TEXT Half Subtractor</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>AA_LABEL</type>
<position>-150.5,-35.5</position>
<gparam>LABEL_TEXT NAND as universal gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>391</ID>
<type>AA_TOGGLE</type>
<position>107.5,-20</position>
<output>
<ID>OUT_0</ID>155 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>392</ID>
<type>AA_TOGGLE</type>
<position>131,-20</position>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_LABEL</type>
<position>-153,-41</position>
<gparam>LABEL_TEXT NAND  as NOT gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>393</ID>
<type>AA_AND2</type>
<position>146,-42</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_AND2</type>
<position>146.5,-52</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>-152.5,-55.5</position>
<gparam>LABEL_TEXT NAND as AND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>396</ID>
<type>AA_INVERTER</type>
<position>115.5,-28</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>203</ID>
<type>BA_NAND2</type>
<position>-159,-65</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>397</ID>
<type>AA_INVERTER</type>
<position>137.5,-27</position>
<input>
<ID>IN_0</ID>156 </input>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>398</ID>
<type>GA_LED</type>
<position>178.5,-45</position>
<input>
<ID>N_in0</ID>162 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>BA_NAND2</type>
<position>-148.5,-65</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>399</ID>
<type>GA_LED</type>
<position>177.5,-56.5</position>
<input>
<ID>N_in0</ID>167 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>400</ID>
<type>AE_OR2</type>
<position>159.5,-44.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>160 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_TOGGLE</type>
<position>-167.5,-64</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>401</ID>
<type>GA_LED</type>
<position>149,-82.5</position>
<input>
<ID>N_in1</ID>166 </input>
<input>
<ID>N_in2</ID>166 </input>
<input>
<ID>N_in3</ID>166 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>402</ID>
<type>GA_LED</type>
<position>149,-91</position>
<input>
<ID>N_in0</ID>165 </input>
<input>
<ID>N_in3</ID>165 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_TOGGLE</type>
<position>-167.5,-67</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>403</ID>
<type>AI_XOR2</type>
<position>143.5,-82.5</position>
<input>
<ID>IN_0</ID>163 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>166 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>GA_LED</type>
<position>-141.5,-65</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>405</ID>
<type>AA_TOGGLE</type>
<position>127,-81</position>
<output>
<ID>OUT_0</ID>163 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>-166.5,-60</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>406</ID>
<type>AA_TOGGLE</type>
<position>124,-83.5</position>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>-167,-70.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>-155,-76</position>
<gparam>LABEL_TEXT NAND as OR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>410</ID>
<type>AA_AND2</type>
<position>145,-60.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>167 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>BA_NAND2</type>
<position>-161.5,-83.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>412</ID>
<type>AA_AND2</type>
<position>143,-91</position>
<input>
<ID>IN_0</ID>168 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>BA_NAND2</type>
<position>-161.5,-90</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>414</ID>
<type>AE_SMALL_INVERTER</type>
<position>135,-90</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_TOGGLE</type>
<position>-168.5,-82.5</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>223</ID>
<type>AA_TOGGLE</type>
<position>-168,-91.5</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>225</ID>
<type>BA_NAND2</type>
<position>-151.5,-86</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>GA_LED</type>
<position>-144,-86</position>
<input>
<ID>N_in0</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>AA_LABEL</type>
<position>-155,-100</position>
<gparam>LABEL_TEXT NAND as NOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>229</ID>
<type>AA_LABEL</type>
<position>-167.5,-78.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>AA_LABEL</type>
<position>-167,-94.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>BA_NAND2</type>
<position>-162,-108</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>233</ID>
<type>BA_NAND2</type>
<position>-162,-114.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>234</ID>
<type>AA_TOGGLE</type>
<position>-169,-107</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>235</ID>
<type>AA_TOGGLE</type>
<position>-168.5,-116</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>236</ID>
<type>BA_NAND2</type>
<position>-152,-110.5</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>BA_NAND2</type>
<position>-142.5,-110.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>GA_LED</type>
<position>-136.5,-110.5</position>
<input>
<ID>N_in2</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>AA_LABEL</type>
<position>-113.5,-43</position>
<gparam>LABEL_TEXT NAND as XOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>BA_NAND2</type>
<position>-108,-49.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>BA_NAND2</type>
<position>-107,-58</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>BA_NAND2</type>
<position>-119.5,-54.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_TOGGLE</type>
<position>-126.5,-48.5</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_TOGGLE</type>
<position>-126,-60.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>254</ID>
<type>BA_NAND2</type>
<position>-99.5,-53</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>256</ID>
<type>GA_LED</type>
<position>-93.5,-53</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>257</ID>
<type>BA_NAND2</type>
<position>-105.5,-78</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>258</ID>
<type>BA_NAND2</type>
<position>-104.5,-86.5</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>259</ID>
<type>BA_NAND2</type>
<position>-117,-83</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>260</ID>
<type>AA_TOGGLE</type>
<position>-124,-77</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_TOGGLE</type>
<position>-123,-89</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>262</ID>
<type>BA_NAND2</type>
<position>-97,-81.5</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>-110.5,-70</position>
<gparam>LABEL_TEXT NAND as XNOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>266</ID>
<type>BA_NAND2</type>
<position>-87.5,-81.5</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>91 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>268</ID>
<type>GA_LED</type>
<position>-81.5,-81.5</position>
<input>
<ID>N_in0</ID>92 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_AND2</type>
<position>-204,-27</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>270</ID>
<type>AA_LABEL</type>
<position>-38.5,-13</position>
<gparam>LABEL_TEXT NOR as universal gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_TOGGLE</type>
<position>-213.5,-26</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>78</ID>
<type>GA_LED</type>
<position>-197.5,-27</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>272</ID>
<type>BE_NOR2</type>
<position>-50.5,-24.5</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_TOGGLE</type>
<position>-213.5,-28</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>-208,-19</position>
<gparam>LABEL_TEXT AND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>274</ID>
<type>GA_LED</type>
<position>-41.5,-24.5</position>
<input>
<ID>N_in3</ID>94 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>-213,-23</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_LABEL</type>
<position>-213.5,-31</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>276</ID>
<type>AA_TOGGLE</type>
<position>-59,-24.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>-190,-26.5</position>
<gparam>LABEL_TEXT Y=A*B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>277</ID>
<type>AA_LABEL</type>
<position>-50.5,-19</position>
<gparam>LABEL_TEXT NOR as NOT gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AE_OR2</type>
<position>-204,-45</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_TOGGLE</type>
<position>-216,-44</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>279</ID>
<type>BE_NOR2</type>
<position>-54.5,-37.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>-216,-46</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>-214,-41</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>281</ID>
<type>BE_NOR2</type>
<position>-44,-37</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>-214,-50</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>-190,-44.5</position>
<gparam>LABEL_TEXT Y=A+B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>283</ID>
<type>AA_TOGGLE</type>
<position>-61.5,-37</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>90</ID>
<type>GA_LED</type>
<position>-198.5,-45</position>
<input>
<ID>N_in3</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>-214,-37</position>
<gparam>LABEL_TEXT OR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>285</ID>
<type>GA_LED</type>
<position>-36.5,-36.5</position>
<input>
<ID>N_in0</ID>97 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_INVERTER</type>
<position>-198,-62</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>286</ID>
<type>AA_LABEL</type>
<position>-50.5,-32</position>
<gparam>LABEL_TEXT NOR as AND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_TOGGLE</type>
<position>-207,-62</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>-188.5,-62</position>
<input>
<ID>N_in0</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>288</ID>
<type>BE_NOR2</type>
<position>-55.5,-50</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>98 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>-215.5,-61.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>-181,-61.5</position>
<gparam>LABEL_TEXT Y=A'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>290</ID>
<type>BE_NOR2</type>
<position>-55,-58.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>-213.5,-57</position>
<gparam>LABEL_TEXT NOT gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>BE_NOR2</type>
<position>-43,-53.5</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>BA_NAND2</type>
<position>-203.5,-76.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>294</ID>
<type>AA_TOGGLE</type>
<position>-64.5,-50</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_TOGGLE</type>
<position>-215.5,-75.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>296</ID>
<type>AA_TOGGLE</type>
<position>-64.5,-60</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>-216,-77.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>298</ID>
<type>GA_LED</type>
<position>-34.5,-53</position>
<input>
<ID>N_in0</ID>102 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>GA_LED</type>
<position>-196,-76</position>
<input>
<ID>N_in0</ID>31 </input>
<input>
<ID>N_in1</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>299</ID>
<type>AA_AND2</type>
<position>-50.5,-75.5</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>-186.5,-77.5</position>
<gparam>LABEL_TEXT Y=A*B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>300</ID>
<type>AA_TOGGLE</type>
<position>-60,-74.5</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>-184,-74</position>
<gparam>LABEL_TEXT ______</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>302</ID>
<type>AA_TOGGLE</type>
<position>-60,-76.5</position>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>303</ID>
<type>AA_LABEL</type>
<position>-59.5,-71.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>-210.5,-68.5</position>
<gparam>LABEL_TEXT NAND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>304</ID>
<type>AA_LABEL</type>
<position>-60,-79.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>-216,-72.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>-216.5,-80.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>307</ID>
<type>BE_NOR2</type>
<position>-41,-75.5</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>BE_NOR2</type>
<position>-202.5,-91</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>309</ID>
<type>GA_LED</type>
<position>-32.5,-74.5</position>
<input>
<ID>N_in0</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_TOGGLE</type>
<position>-212.5,-90</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>310</ID>
<type>AA_LABEL</type>
<position>-48,-67.5</position>
<gparam>LABEL_TEXT NOR as NAND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_TOGGLE</type>
<position>-213,-92</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>312</ID>
<type>BE_NOR2</type>
<position>-60,-94</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>GA_LED</type>
<position>-195.5,-90.5</position>
<input>
<ID>N_in0</ID>34 </input>
<input>
<ID>N_in1</ID>35 </input>
<input>
<ID>N_in3</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>314</ID>
<type>BE_NOR2</type>
<position>-53,-88.5</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>-215,-86</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>-215,-95</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>316</ID>
<type>BE_NOR2</type>
<position>-51.5,-97.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>-186.5,-91.5</position>
<gparam>LABEL_TEXT Y=A+B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_LABEL</type>
<position>-184,-88</position>
<gparam>LABEL_TEXT ______</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>318</ID>
<type>BE_NOR2</type>
<position>-42,-92.5</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>114 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AI_XOR2</type>
<position>-200,-103.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>320</ID>
<type>AA_TOGGLE</type>
<position>-68.5,-89</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_TOGGLE</type>
<position>-211.5,-102.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>322</ID>
<type>AA_TOGGLE</type>
<position>-67.5,-98.5</position>
<output>
<ID>OUT_0</ID>112 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_TOGGLE</type>
<position>-211.5,-104.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>132</ID>
<type>GA_LED</type>
<position>-193,-103.5</position>
<input>
<ID>N_in3</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>326</ID>
<type>BE_NOR2</type>
<position>-34,-93</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>116 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>-181.5,-103.5</position>
<gparam>LABEL_TEXT Y=AB+AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>328</ID>
<type>GA_LED</type>
<position>-27.5,-93</position>
<input>
<ID>N_in1</ID>117 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>329</ID>
<type>AA_LABEL</type>
<position>-57.5,-83</position>
<gparam>LABEL_TEXT NOR as XOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_LABEL</type>
<position>-183.5,-100.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>-175.5,-100.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AO_XNOR2</type>
<position>837,346</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>AO_XNOR2</type>
<position>-139.5,-28</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>337</ID>
<type>BE_NOR2</type>
<position>-58.5,-112</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_TOGGLE</type>
<position>-152,-27</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>338</ID>
<type>BE_NOR2</type>
<position>-50,-107.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>125 </input>
<output>
<ID>OUT</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>339</ID>
<type>BE_NOR2</type>
<position>-50,-115.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_TOGGLE</type>
<position>-152,-29</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>340</ID>
<type>BE_NOR2</type>
<position>-40.5,-110.5</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>AA_TOGGLE</type>
<position>-67,-107</position>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>-133,-28</position>
<input>
<ID>N_in0</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>342</ID>
<type>AA_TOGGLE</type>
<position>-66,-116.5</position>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_LABEL</type>
<position>-120.5,-28.5</position>
<gparam>LABEL_TEXT Y=AB+A'B'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>-162.5,-25.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>-162.5,-28.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_LABEL</type>
<position>-149,-18.5</position>
<gparam>LABEL_TEXT XNOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>346</ID>
<type>GA_LED</type>
<position>-32.5,-110</position>
<input>
<ID>N_in0</ID>131 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>347</ID>
<type>AA_LABEL</type>
<position>-57.5,-102.5</position>
<gparam>LABEL_TEXT NOR as XNOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>349</ID>
<type>AA_LABEL</type>
<position>32.5,-11.5</position>
<gparam>LABEL_TEXT Half Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>355</ID>
<type>AA_TOGGLE</type>
<position>23,-18.5</position>
<output>
<ID>OUT_0</ID>142 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>357</ID>
<type>AA_TOGGLE</type>
<position>46.5,-18.5</position>
<output>
<ID>OUT_0</ID>143 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>359</ID>
<type>AA_AND2</type>
<position>61.5,-40.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>143 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>AA_AND2</type>
<position>62,-50.5</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>363</ID>
<type>AA_AND2</type>
<position>62.5,-59.5</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>143 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>367</ID>
<type>AA_INVERTER</type>
<position>31,-26.5</position>
<input>
<ID>IN_0</ID>142 </input>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_INVERTER</type>
<position>53,-25.5</position>
<input>
<ID>IN_0</ID>143 </input>
<output>
<ID>OUT_0</ID>145 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>371</ID>
<type>GA_LED</type>
<position>94,-43.5</position>
<input>
<ID>N_in0</ID>149 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>373</ID>
<type>GA_LED</type>
<position>93,-55</position>
<input>
<ID>N_in0</ID>148 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>375</ID>
<type>AE_OR2</type>
<position>75,-43</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>377</ID>
<type>AO_XNOR2</type>
<position>-161.5,-37.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>AI_XOR2</type>
<position>44.5,-76.5</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>AA_AND2</type>
<position>45.5,-85</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>BA_NAND2</type>
<position>-150,-47</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>383</ID>
<type>AA_TOGGLE</type>
<position>28,-75</position>
<output>
<ID>OUT_0</ID>150 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_TOGGLE</type>
<position>-162.5,-46</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>385</ID>
<type>AA_TOGGLE</type>
<position>25,-77.5</position>
<output>
<ID>OUT_0</ID>151 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>192</ID>
<type>GA_LED</type>
<position>-141.5,-46.5</position>
<input>
<ID>N_in0</ID>62 </input>
<input>
<ID>N_in1</ID>62 </input>
<input>
<ID>N_in2</ID>62 </input>
<input>
<ID>N_in3</ID>62 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-211.5,-26,-207,-26</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<connection>
<GID>76</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-201,-27,-198.5,-27</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<connection>
<GID>78</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-211.5,-28,-207,-28</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<connection>
<GID>76</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-214,-44,-207,-44</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-214,-46,-207,-46</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-198.5,-45,-198.5,-44</points>
<connection>
<GID>90</GID>
<name>N_in3</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-201,-45,-198.5,-45</points>
<connection>
<GID>84</GID>
<name>OUT</name></connection>
<intersection>-198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-205,-62,-201,-62</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-195,-62,-189.5,-62</points>
<connection>
<GID>94</GID>
<name>N_in0</name></connection>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-213.5,-75.5,-206.5,-75.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-214,-77.5,-206.5,-77.5</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-200.5,-76.5,-195,-76.5</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<intersection>-197 3</intersection>
<intersection>-195 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-197,-76.5,-197,-76</points>
<connection>
<GID>105</GID>
<name>N_in0</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-195,-76.5,-195,-76</points>
<connection>
<GID>105</GID>
<name>N_in1</name></connection>
<intersection>-76.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-210.5,-90,-205.5,-90</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-211,-92,-205.5,-92</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-199.5,-91,-196.5,-91</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>-196.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-196.5,-91,-196.5,-90.5</points>
<connection>
<GID>120</GID>
<name>N_in0</name></connection>
<intersection>-91 1</intersection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-195,-90.5,-195,-89.5</points>
<intersection>-90.5 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-195,-90.5,-194.5,-90.5</points>
<connection>
<GID>120</GID>
<name>N_in1</name></connection>
<intersection>-195 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-195.5,-89.5,-195,-89.5</points>
<connection>
<GID>120</GID>
<name>N_in3</name></connection>
<intersection>-195 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-209.5,-102.5,-203,-102.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-209.5,-104.5,-203,-104.5</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-193,-103.5,-193,-102.5</points>
<connection>
<GID>132</GID>
<name>N_in3</name></connection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-197,-103.5,-193,-103.5</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<intersection>-193 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-150,-27,-142.5,-27</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<connection>
<GID>144</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-150,-29,-142.5,-29</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<connection>
<GID>146</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-136.5,-28,-134,-28</points>
<connection>
<GID>148</GID>
<name>N_in0</name></connection>
<connection>
<GID>142</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-160.5,-46,-153,-46</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-153 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-153,-48,-153,-46</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-141.5,-47.5,-141.5,-45.5</points>
<connection>
<GID>192</GID>
<name>N_in2</name></connection>
<connection>
<GID>192</GID>
<name>N_in3</name></connection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-147,-47,-140.5,-47</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>-142.5 6</intersection>
<intersection>-141.5 0</intersection>
<intersection>-140.5 7</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-142.5,-47,-142.5,-46.5</points>
<connection>
<GID>192</GID>
<name>N_in0</name></connection>
<intersection>-47 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-140.5,-47,-140.5,-46.5</points>
<connection>
<GID>192</GID>
<name>N_in1</name></connection>
<intersection>-47 1</intersection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-153.5,-65,-153.5,-64</points>
<intersection>-65 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-153.5,-64,-151.5,-64</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-153.5 0</intersection>
<intersection>-151.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-156,-65,-153.5,-65</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>-153.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-151.5,-66,-151.5,-64</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>-64 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-145.5,-65,-142.5,-65</points>
<connection>
<GID>211</GID>
<name>N_in0</name></connection>
<connection>
<GID>205</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-165.5,-64,-162,-64</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-163.5,-67,-163.5,-66</points>
<intersection>-67 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-163.5,-66,-162,-66</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>-163.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-165.5,-67,-163.5,-67</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>-163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-166.5,-82.5,-164.5,-82.5</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<connection>
<GID>221</GID>
<name>OUT_0</name></connection>
<intersection>-164.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-164.5,-84.5,-164.5,-82.5</points>
<connection>
<GID>217</GID>
<name>IN_1</name></connection>
<intersection>-82.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-165,-91.5,-165,-91</points>
<intersection>-91.5 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-165,-91,-164.5,-91</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>-165 0</intersection>
<intersection>-164.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-166,-91.5,-165,-91.5</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>-165 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-164.5,-91,-164.5,-89</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>-91 1</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-156.5,-85,-156.5,-83.5</points>
<intersection>-85 1</intersection>
<intersection>-83.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-156.5,-85,-154.5,-85</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>-156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-158.5,-83.5,-156.5,-83.5</points>
<connection>
<GID>217</GID>
<name>OUT</name></connection>
<intersection>-156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-156.5,-90,-156.5,-87</points>
<intersection>-90 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-156.5,-87,-154.5,-87</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>-156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-158.5,-90,-156.5,-90</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<intersection>-156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-148.5,-86,-145,-86</points>
<connection>
<GID>227</GID>
<name>N_in0</name></connection>
<connection>
<GID>225</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-167,-107,-165,-107</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>-165 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-165,-109,-165,-107</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<intersection>-107 1</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-165.5,-116,-165.5,-115.5</points>
<intersection>-116 2</intersection>
<intersection>-115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-165.5,-115.5,-165,-115.5</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<intersection>-165.5 0</intersection>
<intersection>-165 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-166.5,-116,-165.5,-116</points>
<connection>
<GID>235</GID>
<name>OUT_0</name></connection>
<intersection>-165.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-165,-115.5,-165,-113.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>-115.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-157,-109.5,-157,-108</points>
<intersection>-109.5 1</intersection>
<intersection>-108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-157,-109.5,-155,-109.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>-157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-159,-108,-157,-108</points>
<connection>
<GID>232</GID>
<name>OUT</name></connection>
<intersection>-157 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-157,-114.5,-157,-111.5</points>
<intersection>-114.5 2</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-157,-111.5,-155,-111.5</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>-157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-159,-114.5,-157,-114.5</points>
<connection>
<GID>233</GID>
<name>OUT</name></connection>
<intersection>-157 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-147,-111.5,-147,-109.5</points>
<intersection>-111.5 3</intersection>
<intersection>-110.5 2</intersection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-147,-109.5,-145.5,-109.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>-147 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-149,-110.5,-147,-110.5</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<intersection>-147 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-147,-111.5,-145.5,-111.5</points>
<connection>
<GID>239</GID>
<name>IN_1</name></connection>
<intersection>-147 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-136.5,-111.5,-136.5,-110.5</points>
<connection>
<GID>241</GID>
<name>N_in2</name></connection>
<intersection>-110.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-139.5,-110.5,-136.5,-110.5</points>
<connection>
<GID>239</GID>
<name>OUT</name></connection>
<intersection>-136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124.5,-48.5,-111,-48.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<connection>
<GID>250</GID>
<name>OUT_0</name></connection>
<intersection>-122.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-122.5,-53.5,-122.5,-48.5</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>-48.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-117,-60.5,-117,-59</points>
<intersection>-60.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-117,-59,-110,-59</points>
<connection>
<GID>246</GID>
<name>IN_1</name></connection>
<intersection>-117 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-124,-60.5,-117,-60.5</points>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>-122.5 3</intersection>
<intersection>-117 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-122.5,-60.5,-122.5,-55.5</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<intersection>-60.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-110.5,-57,-110.5,-50.5</points>
<intersection>-57 3</intersection>
<intersection>-54.5 2</intersection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-111,-50.5,-110.5,-50.5</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>-110.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-116.5,-54.5,-110.5,-54.5</points>
<connection>
<GID>248</GID>
<name>OUT</name></connection>
<intersection>-110.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-110.5,-57,-110,-57</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>-110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-103.5,-52,-103.5,-49.5</points>
<intersection>-52 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103.5,-52,-102.5,-52</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>-103.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-105,-49.5,-103.5,-49.5</points>
<connection>
<GID>244</GID>
<name>OUT</name></connection>
<intersection>-103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-103,-58,-103,-54</points>
<intersection>-58 2</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,-54,-102.5,-54</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>-103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-104,-58,-103,-58</points>
<connection>
<GID>246</GID>
<name>OUT</name></connection>
<intersection>-103 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-96.5,-53,-94.5,-53</points>
<connection>
<GID>256</GID>
<name>N_in0</name></connection>
<connection>
<GID>254</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-122,-77,-108.5,-77</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>-119.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-119.5,-82,-119.5,-77</points>
<intersection>-82 5</intersection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-120,-82,-119.5,-82</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>-119.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-114.5,-89,-114.5,-87.5</points>
<intersection>-89 2</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-114.5,-87.5,-107.5,-87.5</points>
<connection>
<GID>258</GID>
<name>IN_1</name></connection>
<intersection>-114.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-121,-89,-114.5,-89</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<intersection>-120 3</intersection>
<intersection>-114.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-120,-89,-120,-84</points>
<connection>
<GID>259</GID>
<name>IN_1</name></connection>
<intersection>-89 2</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,-85.5,-108,-79</points>
<intersection>-85.5 3</intersection>
<intersection>-83 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108.5,-79,-108,-79</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-114,-83,-108,-83</points>
<connection>
<GID>259</GID>
<name>OUT</name></connection>
<intersection>-108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-108,-85.5,-107.5,-85.5</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-101,-80.5,-101,-78</points>
<intersection>-80.5 1</intersection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-101,-80.5,-100,-80.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>-101 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-102.5,-78,-101,-78</points>
<connection>
<GID>257</GID>
<name>OUT</name></connection>
<intersection>-101 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-100.5,-86.5,-100.5,-82.5</points>
<intersection>-86.5 2</intersection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-100.5,-82.5,-100,-82.5</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>-100.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-101.5,-86.5,-100.5,-86.5</points>
<connection>
<GID>258</GID>
<name>OUT</name></connection>
<intersection>-100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-94,-81.5,-90.5,-81.5</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<intersection>-90.5 3</intersection>
<intersection>-90.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-90.5,-82.5,-90.5,-80.5</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>-81.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-84.5,-81.5,-82.5,-81.5</points>
<connection>
<GID>268</GID>
<name>N_in0</name></connection>
<connection>
<GID>266</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-25.5,-55,-23.5</points>
<intersection>-25.5 3</intersection>
<intersection>-24.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-23.5,-53.5,-23.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-24.5,-55,-24.5</points>
<connection>
<GID>276</GID>
<name>OUT_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-55,-25.5,-53.5,-25.5</points>
<connection>
<GID>272</GID>
<name>IN_1</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41.5,-24.5,-41.5,-23.5</points>
<connection>
<GID>274</GID>
<name>N_in3</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47.5,-24.5,-41.5,-24.5</points>
<connection>
<GID>272</GID>
<name>OUT</name></connection>
<intersection>-41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58.5,-38.5,-58.5,-36.5</points>
<intersection>-38.5 3</intersection>
<intersection>-37 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58.5,-36.5,-57.5,-36.5</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>-58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-59.5,-37,-58.5,-37</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>-58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-58.5,-38.5,-57.5,-38.5</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>-58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-37.5,-49,-36</points>
<intersection>-37.5 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49,-36,-47,-36</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>-49 0</intersection>
<intersection>-47 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-51.5,-37.5,-49,-37.5</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<intersection>-49 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-47,-38,-47,-36</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<intersection>-36 1</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,-37,-39,-36.5</points>
<intersection>-37 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,-36.5,-37.5,-36.5</points>
<connection>
<GID>285</GID>
<name>N_in0</name></connection>
<intersection>-39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-41,-37,-39,-37</points>
<connection>
<GID>281</GID>
<name>OUT</name></connection>
<intersection>-39 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,-50,-60.5,-49</points>
<intersection>-50 2</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60.5,-49,-58.5,-49</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>-60.5 0</intersection>
<intersection>-58.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-62.5,-50,-60.5,-50</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>-60.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-58.5,-51,-58.5,-49</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<intersection>-49 1</intersection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60,-60,-60,-59.5</points>
<intersection>-60 2</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60,-59.5,-58,-59.5</points>
<connection>
<GID>290</GID>
<name>IN_1</name></connection>
<intersection>-60 0</intersection>
<intersection>-58 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-62.5,-60,-60,-60</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<intersection>-60 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-58,-59.5,-58,-57.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>-59.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-52.5,-49,-50</points>
<intersection>-52.5 1</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49,-52.5,-46,-52.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>-49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-50,-49,-50</points>
<connection>
<GID>288</GID>
<name>OUT</name></connection>
<intersection>-49 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-58.5,-49,-54.5</points>
<intersection>-58.5 2</intersection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49,-54.5,-46,-54.5</points>
<connection>
<GID>292</GID>
<name>IN_1</name></connection>
<intersection>-49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52,-58.5,-49,-58.5</points>
<connection>
<GID>290</GID>
<name>OUT</name></connection>
<intersection>-49 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37.5,-53.5,-37.5,-53</points>
<intersection>-53.5 2</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-37.5,-53,-35.5,-53</points>
<connection>
<GID>298</GID>
<name>N_in0</name></connection>
<intersection>-37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-40,-53.5,-37.5,-53.5</points>
<connection>
<GID>292</GID>
<name>OUT</name></connection>
<intersection>-37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58,-74.5,-53.5,-74.5</points>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58,-76.5,-53.5,-76.5</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<connection>
<GID>299</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45.5,-76.5,-45.5,-74.5</points>
<intersection>-76.5 3</intersection>
<intersection>-75.5 2</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-74.5,-44,-74.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>-45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47.5,-75.5,-45.5,-75.5</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<intersection>-45.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-45.5,-76.5,-44,-76.5</points>
<connection>
<GID>307</GID>
<name>IN_1</name></connection>
<intersection>-45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-75.5,-35.5,-74.5</points>
<intersection>-75.5 2</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,-74.5,-33.5,-74.5</points>
<connection>
<GID>309</GID>
<name>N_in0</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-38,-75.5,-35.5,-75.5</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61,-89,-61,-87.5</points>
<intersection>-89 2</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-61,-87.5,-56,-87.5</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>-61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66.5,-89,-61,-89</points>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection>
<intersection>-63 3</intersection>
<intersection>-61 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-63,-93,-63,-89</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>-89 2</intersection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,-96.5,-55,-89.5</points>
<intersection>-96.5 1</intersection>
<intersection>-94 3</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-96.5,-54.5,-96.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-56,-89.5,-55,-89.5</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-57,-94,-55,-94</points>
<connection>
<GID>312</GID>
<name>OUT</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-65.5,-98.5,-54.5,-98.5</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<connection>
<GID>322</GID>
<name>OUT_0</name></connection>
<intersection>-63 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-63,-98.5,-63,-95</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<intersection>-98.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-47.5,-91.5,-47.5,-88.5</points>
<intersection>-91.5 1</intersection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47.5,-91.5,-45,-91.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>-47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-50,-88.5,-47.5,-88.5</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<intersection>-47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-97.5,-46.5,-93.5</points>
<intersection>-97.5 2</intersection>
<intersection>-93.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46.5,-93.5,-45,-93.5</points>
<connection>
<GID>318</GID>
<name>IN_1</name></connection>
<intersection>-46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-48.5,-97.5,-46.5,-97.5</points>
<connection>
<GID>316</GID>
<name>OUT</name></connection>
<intersection>-46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-94,-38,-92</points>
<intersection>-94 3</intersection>
<intersection>-92.5 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38,-92,-37,-92</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>-38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-39,-92.5,-38,-92.5</points>
<connection>
<GID>318</GID>
<name>OUT</name></connection>
<intersection>-38 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-38,-94,-37,-94</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<intersection>-38 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-31,-93,-26.5,-93</points>
<connection>
<GID>328</GID>
<name>N_in1</name></connection>
<connection>
<GID>326</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,-107,-59.5,-106.5</points>
<intersection>-107 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59.5,-106.5,-53,-106.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>-59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65,-107,-59.5,-107</points>
<connection>
<GID>341</GID>
<name>OUT_0</name></connection>
<intersection>-61.5 3</intersection>
<intersection>-59.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-61.5,-111,-61.5,-107</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>-107 2</intersection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,-114.5,-53.5,-108.5</points>
<intersection>-114.5 1</intersection>
<intersection>-112 3</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-53.5,-114.5,-53,-114.5</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,-108.5,-53,-108.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-55.5,-112,-53.5,-112</points>
<connection>
<GID>337</GID>
<name>OUT</name></connection>
<intersection>-53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,-116.5,-53,-116.5</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<connection>
<GID>339</GID>
<name>IN_1</name></connection>
<intersection>-61.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-61.5,-116.5,-61.5,-113</points>
<connection>
<GID>337</GID>
<name>IN_1</name></connection>
<intersection>-116.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-109.5,-46,-107.5</points>
<intersection>-109.5 1</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46,-109.5,-43.5,-109.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>-46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-107.5,-46,-107.5</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<intersection>-46 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45,-115.5,-45,-111.5</points>
<intersection>-115.5 2</intersection>
<intersection>-111.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45,-111.5,-43.5,-111.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>-45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-115.5,-45,-115.5</points>
<connection>
<GID>339</GID>
<name>OUT</name></connection>
<intersection>-45 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-110.5,-35.5,-110</points>
<intersection>-110.5 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,-110,-33.5,-110</points>
<connection>
<GID>346</GID>
<name>N_in0</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-37.5,-110.5,-35.5,-110.5</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-58.5,23,-20.5</points>
<connection>
<GID>355</GID>
<name>OUT_0</name></connection>
<intersection>-58.5 1</intersection>
<intersection>-49.5 3</intersection>
<intersection>-23.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-58.5,59.5,-58.5</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23,-49.5,59,-49.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>23,-23.5,31,-23.5</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-60.5,46.5,-20.5</points>
<connection>
<GID>357</GID>
<name>OUT_0</name></connection>
<intersection>-60.5 1</intersection>
<intersection>-41.5 2</intersection>
<intersection>-22.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-60.5,59.5,-60.5</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-41.5,58.5,-41.5</points>
<connection>
<GID>359</GID>
<name>IN_1</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>46.5,-22.5,53,-22.5</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-39.5,31,-29.5</points>
<connection>
<GID>367</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-39.5,58.5,-39.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-51.5,53,-28.5</points>
<connection>
<GID>369</GID>
<name>OUT_0</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-51.5,59,-51.5</points>
<connection>
<GID>361</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-42,68,-40.5</points>
<intersection>-42 1</intersection>
<intersection>-40.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-42,72,-42</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-40.5,68,-40.5</points>
<connection>
<GID>359</GID>
<name>OUT</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-50.5,68.5,-44</points>
<intersection>-50.5 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-44,72,-44</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65,-50.5,68.5,-50.5</points>
<connection>
<GID>361</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-59.5,78.5,-55</points>
<intersection>-59.5 2</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-55,92,-55</points>
<connection>
<GID>373</GID>
<name>N_in0</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-59.5,78.5,-59.5</points>
<connection>
<GID>363</GID>
<name>OUT</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-43.5,85.5,-43</points>
<intersection>-43.5 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-43.5,93,-43.5</points>
<connection>
<GID>371</GID>
<name>N_in0</name></connection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-43,85.5,-43</points>
<connection>
<GID>375</GID>
<name>OUT</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-75.5,41.5,-75.5</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>30 10</intersection>
<intersection>33.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>33.5,-84,33.5,-75.5</points>
<intersection>-84 5</intersection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>33.5,-84,42.5,-84</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>33.5 4</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>30,-75.5,30,-75</points>
<connection>
<GID>383</GID>
<name>OUT_0</name></connection>
<intersection>-75.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-86,32,-77.5</points>
<intersection>-86 3</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-77.5,41.5,-77.5</points>
<connection>
<GID>379</GID>
<name>IN_1</name></connection>
<connection>
<GID>385</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32,-86,42.5,-86</points>
<connection>
<GID>381</GID>
<name>IN_1</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-85,50,-85</points>
<connection>
<GID>389</GID>
<name>N_in0</name></connection>
<connection>
<GID>381</GID>
<name>OUT</name></connection>
<intersection>50 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50,-85,50,-84</points>
<connection>
<GID>389</GID>
<name>N_in3</name></connection>
<intersection>-85 1</intersection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-77.5,50,-75.5</points>
<connection>
<GID>387</GID>
<name>N_in3</name></connection>
<connection>
<GID>387</GID>
<name>N_in2</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-76.5,51,-76.5</points>
<connection>
<GID>387</GID>
<name>N_in1</name></connection>
<connection>
<GID>379</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-51,107.5,-22</points>
<connection>
<GID>391</GID>
<name>OUT_0</name></connection>
<intersection>-51 3</intersection>
<intersection>-25 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107.5,-51,143.5,-51</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>107.5,-25,115.5,-25</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-43,131,-22</points>
<connection>
<GID>392</GID>
<name>OUT_0</name></connection>
<intersection>-43 2</intersection>
<intersection>-24 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>131,-43,143,-43</points>
<connection>
<GID>393</GID>
<name>IN_1</name></connection>
<intersection>131 0</intersection>
<intersection>131.5 5</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131,-24,137.5,-24</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>131 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>131.5,-61.5,131.5,-43</points>
<intersection>-61.5 6</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>131.5,-61.5,142,-61.5</points>
<connection>
<GID>410</GID>
<name>IN_1</name></connection>
<intersection>131.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-41,115.5,-31</points>
<connection>
<GID>396</GID>
<name>OUT_0</name></connection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-41,143,-41</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>115 2</intersection>
<intersection>115.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>115,-59.5,115,-41</points>
<intersection>-59.5 3</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>115,-59.5,142,-59.5</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>115 2</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-53,137.5,-30</points>
<connection>
<GID>397</GID>
<name>OUT_0</name></connection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137.5,-53,143.5,-53</points>
<connection>
<GID>394</GID>
<name>IN_1</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,-43.5,152.5,-42</points>
<intersection>-43.5 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152.5,-43.5,156.5,-43.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>152.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>149,-42,152.5,-42</points>
<connection>
<GID>393</GID>
<name>OUT</name></connection>
<intersection>152.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-52,153,-45.5</points>
<intersection>-52 2</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>153,-45.5,156.5,-45.5</points>
<connection>
<GID>400</GID>
<name>IN_1</name></connection>
<intersection>153 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>149.5,-52,153,-52</points>
<connection>
<GID>394</GID>
<name>OUT</name></connection>
<intersection>153 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-45,170,-44.5</points>
<intersection>-45 1</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170,-45,177.5,-45</points>
<connection>
<GID>398</GID>
<name>N_in0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>162.5,-44.5,170,-44.5</points>
<connection>
<GID>400</GID>
<name>OUT</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>129,-81.5,140.5,-81.5</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>129 10</intersection>
<intersection>133 11</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>129,-81.5,129,-81</points>
<connection>
<GID>405</GID>
<name>OUT_0</name></connection>
<intersection>-81.5 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>133,-90,133,-81.5</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<intersection>-81.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126,-83,127.5,-83</points>
<intersection>126 7</intersection>
<intersection>127.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>127.5,-92,127.5,-83</points>
<intersection>-92 8</intersection>
<intersection>-83.5 9</intersection>
<intersection>-83 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>126,-83.5,126,-83</points>
<connection>
<GID>406</GID>
<name>OUT_0</name></connection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>127.5,-92,140,-92</points>
<connection>
<GID>412</GID>
<name>IN_1</name></connection>
<intersection>127.5 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>127.5,-83.5,140.5,-83.5</points>
<connection>
<GID>403</GID>
<name>IN_1</name></connection>
<intersection>127.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,-91,149,-91</points>
<connection>
<GID>412</GID>
<name>OUT</name></connection>
<connection>
<GID>402</GID>
<name>N_in0</name></connection>
<intersection>149 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>149,-91,149,-90</points>
<connection>
<GID>402</GID>
<name>N_in3</name></connection>
<intersection>-91 1</intersection></vsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-83.5,149,-81.5</points>
<connection>
<GID>401</GID>
<name>N_in3</name></connection>
<connection>
<GID>401</GID>
<name>N_in2</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>146.5,-82.5,150,-82.5</points>
<connection>
<GID>403</GID>
<name>OUT</name></connection>
<connection>
<GID>401</GID>
<name>N_in1</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-60.5,162,-56.5</points>
<intersection>-60.5 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162,-56.5,176.5,-56.5</points>
<connection>
<GID>399</GID>
<name>N_in0</name></connection>
<intersection>162 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-60.5,162,-60.5</points>
<connection>
<GID>410</GID>
<name>OUT</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137,-90,140,-90</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<connection>
<GID>414</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>